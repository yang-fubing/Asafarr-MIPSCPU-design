`ifndef __MYCPU_SVH__
`define __MYCPU_SVH__

`include "instr/instr.svh"
`include "cache/cache.svh"
`include "context/context.svh"
`include "mycommon.svh"

`endif
